//U型指令
//LUI
`define LUI_MASK 32'h7F
`define LUI 32'h37
//AUIPC
`define AUIPC_MASK 32'h7F
`define AUIPC 32'h17
//J型指令
//JAL
`define JAL_MASK 32'h7F
`define JAL 32'h6F
//B型指令
//I型指令
//S型指令
//R型指令